/*
 * Copyright (c) 2025 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none


`default_nettype none

// Change the name of this module to something that reflects its functionality and includes your name for uniqueness
// For example tqvp_yourname_spi for an SPI peripheral.
// Then edit tt_wrapper.v line 41 and change tqvp_example to your chosen module name.
module tqvp_adder (
    input         clk,          // Clock - the TinyQV project clock is normally set to 64MHz.
    input         rst_n,        // Reset_n - low to reset.

    input  [7:0]  ui_in,        // The input PMOD, always available.  Note that ui_in[7] is normally used for UART RX.
                                // The inputs are synchronized to the clock, note this will introduce 2 cycles of delay on the inputs.

    output [7:0]  uo_out,       // The output PMOD.  Each wire is only connected if this peripheral is selected.
                                // Note that uo_out[0] is normally used for UART TX.

    input [5:0]   address,      // Address within this peripheral's address space
    input [31:0]  data_in,      // Data in to the peripheral, bottom 8, 16 or all 32 bits are valid on write.

    // Data read and write requests from the TinyQV core.
    input [1:0]   data_write_n, // 11 = no write, 00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    input [1:0]   data_read_n,  // 11 = no read,  00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    
    output [31:0] data_out,     // Data out from the peripheral, bottom 8, 16 or all 32 bits are valid on read when data_ready is high.
    output        data_ready,

    output        user_interrupt  // Dedicated interrupt request for this peripheral
);

    // Implement a 32-bit read/write register at address 0
    reg [31:0] ctrl;
    always @(posedge clk) begin
        if (!rst_n) begin
            ctrl <= 0;
        end else begin
            if (address == 6'h0 ) begin
                if (data_write_n != 2'b11)              ctrl[7:0]   <= data_in[7:0];
                if (data_write_n[1] != data_write_n[0]) ctrl[15:8]  <= data_in[15:8];
                if (data_write_n == 2'b10)              ctrl[31:16] <= data_in[31:16];
            end
        end
    end

    // The bottom 8 bits of the stored data are added to ui_in and output to uo_out.
    reg hsync;
    reg vsync;
    wire visible;
    reg [9:0] pix_x;
    reg [9:0] pix_y;
    
    wire [1:0]R,G,B ;

    wire start = ctrl[0] ;
    
    video_controller u_video_controller(
        .clk      	(clk       ),
        .reset    	(rst_n     ),
        .polarity 	(1'b1      ), // 0 = negative polarity (VGA, SVGA), 1 = positive polarity (XGA, SXGA)
        .hsync    	(hsync     ),
        .vsync    	(vsync     ),
        .visible  	(visible   ),
        .pix_x    	(pix_x     ),
        .pix_y    	(pix_y     )
    );
    

    bg background (
        .clk(clk),
        .rst_n(rst_n),
        .video_active(visible),
        .pix_x(pix_x),
        .pix_y(pix_y),
        .vsync(vsync),
        .R(R),
        .G(G),
        .B(B),
        .start      (start     )
    );


    // Address 0 reads the example data register.  
    // Address 4 reads ui_in
    // All other addresses read 0.
    assign data_out = (address == 6'h0) ? ctrl :
        (address == 6'h4) ? {22'h0,pix_x } :
        (address == 6'h8) ? {22'h0,pix_y } :
        (address == 6'hc) ? {24'h0,uo_out} :
                      32'h0;

    assign uo_out = {vsync, hsync, B, G, R}; 

    // All reads complete in 1 clock
    assign data_ready = 1;
    
    // User interrupt is generated on rising edge of ui_in[6], and cleared by writing a 1 to the low bit of address 8.
    reg example_interrupt;
    reg last_ui_in_6;

    always @(posedge clk) begin
        if (!rst_n) begin
            example_interrupt <= 0;
        end

        if (ui_in[6] && !last_ui_in_6) begin
            example_interrupt <= 1;
        end else if (address == 6'h8 && data_write_n != 2'b11 && data_in[0]) begin
            example_interrupt <= 0;
        end

        last_ui_in_6 <= ui_in[6];
    end

    assign user_interrupt = example_interrupt;

    // List all unused inputs to prevent warnings
    // data_read_n is unused as none of our behaviour depends on whether
    // registers are being read.
    wire _unused = &{data_read_n, 1'b0};

endmodule

